class tb_sequencer extends uvm_sequencer#(my_trans);

    `uvm_component_utils(tb_sequencer)

    function new (string name = "tb_sequencer",uvm_component parent);
        super.new(name,parent);
    endfunction

endclass

