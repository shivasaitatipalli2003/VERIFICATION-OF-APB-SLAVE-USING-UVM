`include "uvm_macros.svh"

package apb_pkg;

    import uvm_pkg::*;

    `include "apb_uvm_transaction.sv"
    `include "apb_uvm_sequence.sv"
    `include "apb_uvm_sequencer.sv"
    `include "apb_uvm_driver.sv"
    `include "apb_uvm_monitor.sv"
    `include "apb_uvm_prd.sv"
    `include "apb_uvm_cmp.sv"
    `include "apb_uvm_scoreboard.sv"
    `include "apb_uvm_agent.sv"
    `include "apb_uvm_environment.sv"
    `include "apb_uvm_base_test.sv"

endpackage

